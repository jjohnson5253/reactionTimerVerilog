//Jake Johnson 2016

//Reaction timer circuit made for ECEN 2350: Digital Logic

//This reactionTimer is a finite state machine with 3 states
//State 1 (Q=1): LED OFF, NO Timer counting
	//default state
//State 2 (Q=2): LED off, Random generator timer counting, No timer counting
	//reaction timer started, once random time counted the machine will enter state 3
//State 3 (Q-3): LED ON, timer counting
	//LED on and time counts until user presses button to go back to state 1

module reactionTimer(Clock, Reset, Pushn, LED, LED2, LED3, LED4,LED5, Digit1, Digit0);

	input Clock, Reset,Pushn;
	output reg LED, LED2, LED5;
	output LED3, LED4;

	output wire [1:7]Digit1,Digit0;	//sev seg display values				
	wire [3:0]BCD1,BCD0; //counter number					
	wire c9; 		//divided clock signal					
	reg[1:0]Q = 1;	//state variable	
	wire [3:0]randomNumber;	 //random number generated by LFSR	
	reg enableCount, enableLFSR;
	wire doneCount;
	reg lastPush;
	reg ss;
	wire [10:0]mycounter;
	initial lastPush = ss;
	wire [10:0] val;
	assign val = 150;

	always@(posedge !Pushn) //change state of button pressed variable 'ss'
	begin
		ss = !ss;
	end
	
	always@(posedge Clock)
	begin
	
		if(ss!=lastPush) //if button variable is different then before it was pushed..
		begin
			case(Q)
			1 : Q <= 2;
			2 : ;
			3 : Q <= 1;
			endcase
			lastPush=ss;
		end
		/*
		if(doneCount)begin
			if(Q==2)begin
				LED5<=1;
			end
		end*/

		case(Q)
		1: begin
			LED<=0; //LED OFF (LED CONTROLS IF LIGHT IS ON AND IF COUNTER IS ENABLED)
			LED2<=0;
			enableLFSR <= 1;
			enableCount <= 0;
			end
		2: begin
			LED<=0; //LED OFF
			//LED2<=1;
			enableLFSR <= 0;
			enableCount <= 1;
			if(doneCount) begin
				Q <= 3;
				LED5<=0;
			end
			else
				LED5<=0;
			end
		3: begin
			LED<=1; //LED ON
			LED2<=0;
			enableLFSR<=0;
			enableCount<=0;
			end
		endcase
	
	end
	
	clockDivider hundredHertz(Clock,c9); //divide clock to get our frequency
	BCDcount counter(c9,Reset,LED,BCD1,BCD0,LED4);
	seg7 seg1(BCD1,Digit1);
	seg7 seg0(BCD0,Digit0);

	//LFSR ranNum(Clock,enableLFSR,randomNumber, LED4);
	countTo count1(c9, val, doneCount, enableCount, LED3, mycounter);

endmodule

//////////////////////////////////////////////////////////////////////////////

module BCDcount(Clock,Clear,E,BCD1,BCD0,LED4);
	input Clock,Clear,E;
	output reg [3:0]BCD1,BCD0;
	output reg LED4;
	initial LED4 = 0;
	always@(posedge Clock)
	begin
		if(Clear) //if clear, set everything to 0
		begin
			BCD1<=0;
			BCD0<=0;
		end
		else if(~Clear && E) //if enable... NOTE: this module is enabled by the LED
			if(BCD0==4'b1001)//if BCD0 is 9 (right digit)
			begin
				BCD0<=0; //set it back to 0
				if(BCD1==4'b1001) //if BCD1 9
					BCD1<=0; //set back to 0
				else 
					BCD1<=BCD1+1; //otherwise increment
			end
		else 
			BCD0<=BCD0+1; //if !Clear and E, then increment BCD0
	end

	//note: as long as BCD0!=9, it increments on clockedge 
	//and BCD1 remains in its state, so BCDO goes up to 9
	//before BCD1 increments


	//ALSO: I think we could just add another BCD (BCD2) and make that 
	//increment everytime BCD1 gets to 9 (just put this incrementation 
	//inside an if statement exactly like what we did for BCD1 and BCD0)

endmodule

/////////////////////////////////////////////////////////////////////////

module seg7(bcd,leds);
	input [3:0]bcd;
	output reg[1:7] leds;

	always@(bcd)
		case(bcd)  //whenever bcd changes, change led outputs accordingly
					  //abcdefg
			0: leds=7'b0000001;//1111110;
			1: leds=7'b1001111;//0110000;
			2: leds=7'b0010010;//1101101;
			3: leds=7'b0000110;//1111001;
			4: leds=7'b1001100;//0110011;
			5: leds=7'b0100100;//1011011;
			6: leds=7'b0100000;//1011111;
			7: leds=7'b0001111;//1110000;
			8: leds=7'b0000000;//1111111;
			9: leds=7'b0000100;//1111011;
			default: leds=7'bx;
		endcase

endmodule


//////////////////////Clock Divider///////////////////////////////////////////////////////
////////////takes in Clock and effectively outputs that frequency%10 ///////////////////////


module clockDivider(Clock,c19);
	input Clock;
	reg [19:0]Q;
	output reg c19;

	always@(posedge Clock)
	begin
		Q <= Q+1;
		
		c19 = Q[19];
	end

endmodule

////////////////////////////////////////////////////////////////////////////
/*
//this linear feedback shift register will produce a psuedo random number
module LFSR(Clock,enable,num,LED);
input Clock,enable;
output reg [3:0] num;
output reg LED;
initial num = 1;

always@(posedge Clock)
begin
	if(enable)
	begin
		LED = 1;
		num[3] = num[3] ^ num[0];
		num[2] = num[3];
		num[1] = num[2];
		num[0] = num[1];
	end
	else
		LED = 0;
end
endmodule
*/
///////////////////////////////////////////////////////////////////////////////

module countTo(clock, inputN, done, enable, LED3, counter);
	input clock, enable;
	input [10:0] inputN;
	output reg done;
	output reg LED3;
	output reg[10:0]counter;
	initial counter = 1;
	initial LED3 = 0;
	initial done = 0;
	//reg [10:0] test;
	//initial test = 20;
	//wire [10:0] test;
	//assign test = inputN;
	
	always@(posedge clock)
	begin
	
		if(enable)
		begin
			case(counter)
			inputN : begin
				done <= 1;
				//LED3 <= 1;
				end
			200 : begin
				counter = 1;
				end
			default : begin
				counter<=counter+1;
				LED3<=0;
				end
			endcase
		end
		else begin
			LED3 <= 0;
		end
	end
endmodule








